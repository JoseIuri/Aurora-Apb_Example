package arith_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    

    `include "apb_coverage.sv"
	`include "apb_driver.sv"
	`include "apbSequence_sequence.sv"
	`include "apb_transaction.sv"
	`include "arith_scoreboard.sv"
	`include "apbTest_test.sv"
	`include "arith_env.sv"
	`include "arithRefmod_refmod.sv"
	`include "apb_agent.sv"
	`include "apb_monitor.sv"
	
endpackage